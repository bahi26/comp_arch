library ieee;
use ieee.std_logic_1164.all;
entity forward_unit is
	port(mem_input,wb_input:in std_logic_vector(5 downto 0);
	     s13_mem,s13_wb:in std_logic_vector(1 downto 0);
	     rs,rd:in std_logic_vector(2 downto 0);
	     esp,msp,wsp:in std_logic;
	     f1,f2:out std_logic_vector(2 downto 0));
end entity forward_unit;
architecture forward_unit_arch of forward_unit is
begin
	f2<="110"  when(esp=msp and esp='1')
	else "111" when(esp=wsp and esp='1')
	else "001" when(mem_input(5 downto 3)=rs and s13_mem(1)='1')
	else "100" when(mem_input(2 downto 0)=rs and s13_mem(0)='1')
	else "011" when(wb_input(5 downto 3)=rs and s13_wb(1)='1')
	else "101" when(wb_input(2 downto 0)=rs and s13_wb(0)='1')
	else "000";
	f1<= "001" when(mem_input(5 downto 3)=rd and s13_mem(1)='1')
	else "100" when(mem_input(2 downto 0)=rd and s13_mem(0)='1')
	else "011" when(wb_input(5 downto 3)=rd and s13_wb(1)='1')
	else "101" when(wb_input(2 downto 0)=rd and s13_wb(0)='1')
	else "000";
end forward_unit_arch;